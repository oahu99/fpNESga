module color_palette
(
    input logic [7:0] palette_address,
    output logic [7:0] r, g, b
);